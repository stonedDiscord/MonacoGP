.title KiCad schematic
.include "/home/stoned/MonacoGP/7400.LIB"
.include "/home/stoned/MonacoGP/IC.LIB"
.model __D3 D
.model __D1 D
.model __D2 D
.model __Q1 NPN level=4
.save all
.probe alli
XU58 _BRIDGE_AP _M-ROAD Net-_U58-Pad3_ 7408
XU72 Net-_U117-Pad1_ Net-_U119-Za_ _WALL 7400
XU97 7442
XU98 MH0 Net-_U98-I0a_ Net-_U98-I1a_ Net-_U97-A0_ Net-_U98-I0b_ Net-_U98-I1b_ Net-_U97-A1_ GNDPWR Net-_U97-A2_ Net-_U98-I1c_ Net-_U98-I0c_ unconnected-_U98-Zd-Pad12_ Net-_U98-I1d_ Net-_U98-I0d_ VCC VCC NC-U98-0 NC-U98-1 NC-U98-2 NC-U98-3 NC-U98-4 NC-U98-5 NC-U98-6 74157
XU119 74153
XU120 EPROM_2716
XU99 EPROM_2716
XU48 VCC VCC _MHL0 Net-_U40B-D_ Net-_U48-Z_ unconnected-_U48-_Z-Pad6_ GNDPWR GNDPWR Net-_U41-S2_ Net-_U41-S1_ Net-_U41-S0_ Net-_U40B-D_ VCC VCC VCC 74151
XU40 Net-_U25A-_R_ EXTEND Net-_U24-0_ unconnected-_U40A-_S-Pad4_ Net-_U40A-Q_ Net-_U40A-_Q_ 7474
XU74 _M2VL0 FN _M1VL0 unconnected-_U74A-_S-Pad4_ E7 _ROAD 7474
C1 _ROAD GNDPWR 470p
XU45 Net-_U40B-_Q_ Net-_U38A-Q_ Net-_U25B-_R_ 7400
XU86 AREA_5 unconnected-_U86-I6-Pad14_ Net-_U79-D2_ GNDPWR VCC 74368
XU80 BRIDGE_AP Net-_U25A-_Q_ Net-_U68B-Q_ 7402
XU117 Net-_U117-Pad1_ Net-_U120-A8_ 7406
XU87 EA Net-_U87-Pad2_ Net-_U83-S_ 7408
XU89 7427
XU104 EN Net-_U88B-Q_ Net-_U67-S_ 7432
XU204 Net-_U204-Pad1_ Net-_U204-Pad2_ Net-_U202-I0d_ 7486
C25 Net-_U202-I0d_ GNDPWR 470p
XU55 _DUMMY__W_ Net-_U52-Pad10_ E6 FF 7410
XU90 M2V1 M2V0 NC-U90-0 Net-_U117-Pad4_ M2V4 7420
XU81 Net-_U81-Pad1_ Net-_U81-Pad2_ FC 7400
XU88 Net-_U88A-_R_ MH6 MH5 unconnected-_U88A-_S-Pad4_ unconnected-_U88A-Q-Pad5_ Net-_U88A-_Q_ 7474
XU82 Net-_U78-Pad8_ Net-_U81-Pad1_ 7406
XU201 74393
XU78 M1V0 M1V1 NC-U78-0 M1V4 M1V3 7420
XU59 EM Net-_U46-DOWN_ 7406
XU94 EW E20 Net-_U96-0_ _Y-LINE 7410
XU73 7427
XU202 Net-_U201A-MR_ Net-_U201B-Q0_ D17 S-100-A Net-_U201B-Q1_ D16 S-100-B GNDPWR S-100-D D15 Net-_U201B-Q2_ S-100-C D14 Net-_U202-I0d_ VCC VCC NC-U202-0 NC-U202-1 NC-U202-2 NC-U202-3 NC-U202-4 NC-U202-5 NC-U202-6 74157
RN1 VCC D10 560
XU205 Net-_U201A-MR_ GNDPWR F16 SP.A GNDPWR FT SP.B GNDPWR SP.C F17 GNDPWR SP.D FU Net-_U205-I0d_ VCC VCC NC-U205-0 NC-U205-1 NC-U205-2 NC-U205-3 NC-U205-4 NC-U205-5 NC-U205-6 74157
XU101 FF GNDPWR NC-U101-0 Net-_U107-D0_ Net-_U101-Pad5_ 7420
XU203 Net-_U201A-MR_ Net-_U201B-Q3_ EB EXTEND Net-_U203-I0b_ E3 _EXTEND GNDPWR ED E6 Net-_U201A-MR_ unconnected-_U203-Zd-Pad12_ unconnected-_U203-I1d-Pad13_ unconnected-_U203-I0d-Pad14_ VCC VCC NC-U203-0 NC-U203-1 NC-U203-2 NC-U203-3 NC-U203-4 NC-U203-5 NC-U203-6 74157
XU206 ED Net-_U206A-D_ F19 unconnected-_U206A-_S-Pad4_ unconnected-_U206A-Q-Pad5_ Net-_U206A-D_ 7474
XU46 74193
XU39 unconnected-_U39-Pad1_ unconnected-_U39-Pad2_ unconnected-_U39-Pad3_ 7432
XU52 Net-_U46-QB_ Net-_U46-QA_ Net-_U39-Pad4_ 7408
C5 _DUMMY_AREA GNDPWR 470p
XU56 Net-_U68B-Q_ Net-_U104-Pad11_ Net-_U56-Pad12_ 7400
XU42 FG F7 V-CA Vb 7410
XU65 Net-_U65-Pad1_ EJ V-4 7402
XU26 _SIG.__BL_ _DUMMY__BL_ NC-U26-0 EU Net-_U19-Pad6_ 7420
XU60 7427
XU61 7427
XU47 VCC FJ Net-_U40B-D_ 7408
XU49 74393
XU62 Net-_U61-Pad6_ Net-_U69B-_R_ 7406
XU93 E21 _V4 7406
XU53 74153
XU66 _DUMMY_AREA E9 Net-_U66-Pad3_ _0-AREA 7410
XU9 Net-_U50-Zd_ Net-_U66-Pad8_ _SIG.__Y_ 7400
XU16 Net-_U16-Pad1_ Net-_U15-Pad8_ F4 7400
XU50 H0 Net-_U50-I0a_ Net-_U50-I1a_ Net-_U50-Za_ Net-_U50-I0b_ Net-_U50-I1b_ Net-_U50-Zb_ GNDPWR unconnected-_U50-Zc-Pad9_ Net-_U50-I1c_ Net-_U50-I0c_ Net-_U50-Zd_ Net-_U50-I1d_ Net-_U50-I0d_ VCC VCC NC-U50-0 NC-U50-1 NC-U50-2 NC-U50-3 NC-U50-4 NC-U50-5 NC-U50-6 74157
XU51 EPROM_2716
XU115 V2 FF _H5 FG 7410
XU116 Net-_U107-D1_ FB FF Net-_U107-D0_ Net-_U107-D0_ Net-_U107-D1_ FF FF 74107
XU114 FF FN 7406
XU41 Net-_U40B-D_ Net-_U40B-D_ Net-_U40B-D_ VCC Net-_U41-Z_ unconnected-_U41-_Z-Pad6_ GNDPWR GNDPWR Net-_U41-S2_ Net-_U41-S1_ Net-_U41-S0_ _MHL0 Net-_U40B-D_ Net-_U40B-D_ VCC 74151
C2 V-CA GNDPWR 470p
C13 Net-_U100-_PE_ GNDPWR 470p
XU100 VCC Net-_U100-CP_ Net-_U100-D0_ Net-_U100-D0_ Net-_U100-D0_ Net-_U100-D0_ VCC GNDPWR Net-_U100-_PE_ Net-_U100-CET_ EN E12 V5 E21 V-CA VCC NC-U100-0 NC-U100-1 NC-U100-2 74161
XU110 V-CA FF FS 7400
XU28 Net-_U16-Pad1_ E21 Net-_U21-Pad11_ 7486
C8 F12 GNDPWR 470p
C19 Net-_U100-CP_ GNDPWR 470p
XU1 Net-_U1-Pad1_ Net-_R6-Pad1_ 7407
XU109 VCC Net-_U100-D0_ FF VCC Net-_U109B-Q_ 7MHz VCC VCC 74107
C998 V-CA GNDPWR 470p
XU102 VCC Net-_U100-CP_ GNDPWR GNDPWR GNDPWR FF VCC GNDPWR Net-_U100-_PE_ VCC V3 V2 V1 V0 VCC VCC NC-U102-0 NC-U102-1 NC-U102-2 74161
XU107 VCC 7MHz Net-_U107-D0_ Net-_U107-D1_ GNDPWR VCC Net-_U107-CEP_ GNDPWR Net-_U107-_PE_ VCC H7 FG F7 F8 VCC VCC NC-U107-0 NC-U107-1 NC-U107-2 74161
XU95 VCC Net-_U100-CP_ FJ 7408
Cp19 GNDPWR VCC 100n
Cp24 GNDPWR VCC 100n
Cp20 GNDPWR VCC 100n
Cp21 GNDPWR VCC 100n
Cp26 GNDPWR VCC 100n
Cp33 GNDPWR VCC 100n
Cp32 GNDPWR VCC 100n
Cp28 GNDPWR VCC 100n
Cp30 GNDPWR VCC 100n
Cp31 GNDPWR VCC 100n
Cp25 GNDPWR VCC 100n
Cp34 GNDPWR VCC 100n
Cp23 GNDPWR VCC 100n
Cp29 GNDPWR VCC 100n
Cp27 GNDPWR VCC 100n
Cp22 GNDPWR VCC 100n
Cp36 GNDPWR VCC 100n
Cp35 GNDPWR VCC 100n
J1 __J1
J3 __J3
J2 __J2
XU18 unconnected-_U18A-A-Pad1_ unconnected-_U18A-B-Pad2_ unconnected-_U18A-Clr-Pad3_ unconnected-_U18A-_Q-Pad4_ Net-_U18B-Q_ Net-_U18B-Cext_ Net-_U18B-RCext_ Net-_U18B-A_ Net-_U18B-A_ 74123
XU8 E15 Net-_U19-Pad5_ Net-_U20-Za_ unconnected-_U8-Pad4_ 7410
XU23 V3 Net-_U16-Pad1_ Net-_U12-A3_ 7486
XU3 Net-_U26-Pad6_ Net-_U2-E8_ 7404
Cp7 GNDPWR VCC 100n
Cp14 GNDPWR VCC 100n
Cp11 GNDPWR VCC 100n
Cp12 GNDPWR VCC 100n
Cp1 GNDPWR VCC 100n
Cp2 GNDPWR VCC 100n
Cp13 GNDPWR VCC 100n
Cp9 GNDPWR VCC 100n
Cp15 GNDPWR VCC 100n
Cp6 GNDPWR VCC 100n
Cp10 GNDPWR VCC 100n
Cp5 GNDPWR VCC 100n
Cp8 GNDPWR VCC 100n
Cp4 GNDPWR VCC 100n
Cp3 GNDPWR VCC 100n
Cp16 GNDPWR VCC 100n
Cp18 GNDPWR VCC 100n
Cp17 GNDPWR VCC 100n
XU19 Net-_U10-Pad8_ Net-_U79-Q0_ EC TUNNEL_AP 7410
XU21 V-4 _DUMMY_AREA _HOUSE_ST _GRASSAREA 7411
XU7 _TV-BLANKING Net-_Q1-B_ 7406
XU22 V-4 Net-_U11-E_ 7406
XU15 _ROAD EC Net-_U10-Pad2_ 7408
XU4 E8 unconnected-_U4-Pad2_ Net-_U20-Zd_ unconnected-_U4-Pad4_ E4 Net-_U79-Q3_ GNDPWR Net-_U3-Pad5_ NC-U4-0 7430
XU14 Net-_U14-Pad1_ Net-_U5-Za_ NC-U14-0 7MHz Net-_U13-Pad3_ 7420
XU44 _BRIDGE__R_ _WALL Net-_U57B-Q_ Net-_U37-Q2_ 7410
XU32 7421
XU10 Net-_U10-Pad1_ Net-_U10-Pad2_ Net-_U20-I0b_ 7432
XU31 Net-_U25A-_R_ Net-_U31A-D_ Net-_U24-2_ unconnected-_U31A-_S-Pad4_ Net-_U31A-Q_ Net-_U31A-_Q_ 7474
XU27 _DUMMY__W_ _RESCUE__W_ Net-_U5-Zd_ unconnected-_U27-Pad4_ E17 Net-_U20-Zb_ GNDPWR Net-_U27-Pad8_ NC-U27-0 7430
XU33 _RESCUE__R_ _DUMMY__R_ unconnected-_U33-Pad3_ Net-_TP1-Pad1_ EK ET GNDPWR Net-_U3-Pad11_ NC-U33-0 7430
XU34 Net-_U3-Pad13_ EXTEND Net-_U20-I0b_ 7402
XU25 Net-_U25A-_R_ EXT._500 F3 unconnected-_U25A-_S-Pad4_ Net-_U25A-Q_ Net-_U25A-_Q_ 7474
XU13 unconnected-_U13-Pad1_ _TREE&GRASS__BL_ Net-_U13-Pad3_ _Y-LINE Net-_U2-E9_ Net-_U2-E6_ GNDPWR Net-_U10-Pad1_ NC-U13-0 7430
XU24 7442
C17 Net-_C17-Pad1_ Net-_C17-Pad2_ 0.1u
C16 Net-_C16-Pad1_ Net-_C16-Pad2_ 100p
Y1 __Y1
R18 Net-_C17-Pad2_ Net-_C16-Pad2_ 330
R17 Net-_R17-Pad1_ Net-_C17-Pad1_ 330
XU57 VCC unconnected-_U57A-_Q-Pad2_ MH8 VCC Net-_U57B-Q_ unconnected-_U57B-_Q-Pad6_ VCC VCC 74107
XU35 unconnected-_U35A-_R-Pad1_ FJ Net-_U35A-C_ Net-_U35A-_S_ Net-_U35A-Q_ Net-_U35A-_Q_ 7474
XU38 unconnected-_U38A-_R-Pad1_ Net-_U38A-D_ Net-_U201A-CP_ unconnected-_U38A-_S-Pad4_ Net-_U38A-Q_ Net-_U31A-D_ 7474
R2077 14MHz_EXT VCC 470
XU108 VCC 7MHz GNDPWR GNDPWR GNDPWR Net-_U107-D0_ VCC GNDPWR Net-_U107-_PE_ VCC H3 H2 H1 H0 VCC VCC NC-U108-0 NC-U108-1 NC-U108-2 74161
C14 Net-_U107-_PE_ GNDPWR 470p
XU2 Net-_U2-E4_ Net-_U2-E5_ Net-_U2-E6_ Net-_U2-E7_ Net-_U2-E8_ Net-_U2-S2_ Net-_U2-S1_ GNDPWR Net-_U2-S0_ Net-_U2-E9_ unconnected-_U2-E1-Pad11_ Net-_U2-E2_ Net-_U2-E3_ unconnected-_U2-S3-Pad14_ NC-U2-0 VCC NC-U2-1 74147
R3 VCC D12 470
R1 VCC D11 470
XU79 74174
XU20 EXTEND _TREE&GRASS__G_ unconnected-_U20-I1a-Pad3_ Net-_U20-Za_ Net-_U20-I0b_ _TREE&GRASS__G_ Net-_U20-Zb_ GNDPWR Net-_U20-Zc_ Net-_U20-I1c_ _GRASS Net-_U20-Zd_ _TREE&GRASS__BL_ Net-_U20-I0d_ VCC VCC NC-U20-0 NC-U20-1 NC-U20-2 NC-U20-3 NC-U20-4 NC-U20-5 NC-U20-6 74157
R6 Net-_R6-Pad1_ D13 470
R4 Net-_R4-Pad1_ D12 470
R2 Net-_R2-Pad1_ D11 470
R5 VCC D13 470
D3 D13 Net-_D1-K_ __D3
R13 GNDPWR D11 10k
R14 GNDPWR D12 10k
R15 GNDPWR D13 10k
D1 D11 Net-_D1-K_ __D1
D2 D12 Net-_D1-K_ __D2
Q1 GNDPWR Net-_D1-K_ Net-_Q1-B_ __Q1
XU112 74153
XU113 EPROM_2716
XU43 Net-_U43-S_ GNDPWR GNDPWR Net-_U36-D0_ VCC GNDPWR Net-_U36-D1_ GNDPWR Net-_U36-D2_ GNDPWR GNDPWR Net-_U36-D3_ VCC VCC VCC VCC NC-U43-0 NC-U43-1 NC-U43-2 NC-U43-3 NC-U43-4 NC-U43-5 NC-U43-6 74157
C9 Net-_U43-S_ GNDPWR 470p
R16 Net-_U18B-RCext_ VCC 47k
C4 Net-_U18B-RCext_ Net-_U18B-Cext_ 1.5u
XU30 EPROM_2716
XU105 74153
XU106 EPROM_2716
XU37 VCC 7MHz VCC VCC GNDPWR GNDPWR VCC GNDPWR Net-_U36-_PE_ Net-_U36-TC_ Net-_U37-Q3_ Net-_U37-Q2_ Net-_U30-A7_ Net-_U30-A6_ VCC VCC NC-U37-0 NC-U37-1 NC-U37-2 74161
C6 Net-_U35A-_S_ GNDPWR 470p
XU68 unconnected-_U68A-_R-Pad1_ unconnected-_U68A-_S1-Pad2_ unconnected-_U68A-_S2-Pad3_ unconnected-_U68A-Q-Pad4_ Net-_U41-Z_ Net-_U48-Z_ Net-_U68B-Q_ 74279
XU54 7442
XU69 Net-_U69A-_R_ unconnected-_U69A-D-Pad2_ unconnected-_U69A-C-Pad3_ Net-_U69A-_S_ Net-_U69A-Q_ Net-_U69A-_Q_ 7474
C22 Net-_U54-6_ GNDPWR 470p
XU83 Net-_U83-S_ VCC GNDPWR Net-_U83-Za_ Net-_U69B-Q_ GNDPWR Net-_U83-Zb_ GNDPWR Net-_U83-Zc_ GNDPWR Net-_U69B-Q_ Net-_U83-Zd_ VCC Net-_U69B-_Q_ VCC VCC NC-U83-0 NC-U83-1 NC-U83-2 NC-U83-3 NC-U83-4 NC-U83-5 NC-U83-6 74157
XU29 Net-_U29-S_ Net-_U29-I0a_ Net-_U29-I1a_ Net-_U29-Za_ Net-_U29-I0b_ Net-_U29-I1b_ Net-_U29-Zb_ GNDPWR Net-_U29-Zc_ Net-_U29-I1c_ Net-_U29-I0c_ Net-_U29-Zd_ Net-_U29-I1d_ Net-_U29-I0d_ VCC VCC NC-U29-0 NC-U29-1 NC-U29-2 NC-U29-3 NC-U29-4 NC-U29-5 NC-U29-6 74157
XU84 Net-_U83-S_ VCC GNDPWR Net-_U84-Za_ Net-_U69A-Q_ GNDPWR Net-_U84-Zb_ GNDPWR Net-_U84-Zc_ GNDPWR Net-_U69A-Q_ Net-_U84-Zd_ VCC Net-_U69A-_Q_ VCC VCC NC-U84-0 NC-U84-1 NC-U84-2 NC-U84-3 NC-U84-4 NC-U84-5 NC-U84-6 74157
C12 _M1VL0 GNDPWR 470p
XU70 _M2VL0 V-5 Net-_U69A-_S_ 7432
C7 Net-_U35A-C_ GNDPWR 470p
C18 GNDPWR Net-_U36-_PE_ 470p
XU36 VCC 7MHz Net-_U36-D0_ Net-_U36-D1_ Net-_U36-D2_ Net-_U36-D3_ VCC GNDPWR Net-_U36-_PE_ VCC Net-_U30-A5_ Net-_U30-A4_ Net-_U29-S_ unconnected-_U36-Q0-Pad14_ VCC VCC NC-U36-0 NC-U36-1 NC-U36-2 74161
XU6 7442
XU11 MH0 Net-_U11-I0a_ Net-_U11-I1a_ Net-_U11-Za_ Net-_U11-I0b_ Net-_U11-I1b_ Net-_U11-Zb_ GNDPWR Net-_U11-Zc_ Net-_U11-I1c_ Net-_U11-I0c_ unconnected-_U11-Zd-Pad12_ Net-_U11-I1d_ Net-_U11-I0d_ VCC VCC NC-U11-0 NC-U11-1 NC-U11-2 NC-U11-3 NC-U11-4 NC-U11-5 NC-U11-6 74157
XU12 EPROM_2716
XU17 EPROM_2716
C333 Net-_C333-Pad1_ GNDPWR 470p
XU5 BRIDGE_AP E7 Net-_U5-I1a_ Net-_U5-Za_ E7 _BRIDGE__Bu_ Net-_U5-Zb_ GNDPWR Net-_U5-Zc_ _BRIDGE__Y_ _Y-LINE Net-_U5-Zd_ EG _SIDE_LINE GNDPWR VCC NC-U5-0 NC-U5-1 NC-U5-2 NC-U5-3 NC-U5-4 NC-U5-5 NC-U5-6 74157
XU92 Net-_U67-S_ M1V0 M2V0 Net-_U106-A0_ M1V1 M2V1 Net-_U106-A1_ GNDPWR Net-_U106-A2_ M2V2 M1V2 Net-_U106-A3_ M2V3 M1V3 VCC VCC NC-U92-0 NC-U92-1 NC-U92-2 NC-U92-3 NC-U92-4 NC-U92-5 NC-U92-6 74157
XU67 Net-_U67-S_ M1V4 M2V4 Net-_U106-A4_ _M1VL0 _M2VL0 Net-_U67-Zb_ GNDPWR unconnected-_U67-Zc-Pad9_ unconnected-_U67-I1c-Pad10_ unconnected-_U67-I0c-Pad11_ unconnected-_U67-Zd-Pad12_ unconnected-_U67-I1d-Pad13_ unconnected-_U67-I0d-Pad14_ VCC VCC NC-U67-0 NC-U67-1 NC-U67-2 NC-U67-3 NC-U67-4 NC-U67-5 NC-U67-6 74157
C24 Net-_U40B-_Q_ GNDPWR 470p
C20 ED GNDPWR 470p
XU75 unconnected-_U75-Pad1_ unconnected-_U75-Pad2_ M2V6 M2V7 7410
XU96 7442
TP1 __TP1
XU71 F8 H7 NC-U71-0 FG Net-_U68D-Q_ 7420
XU63 Net-_U63-I3_ Net-_U63-I2_ Net-_U63-I1_ Net-_U63-I0_ unconnected-_U63-Z-Pad5_ Net-_U63-_Z_ Net-_U63-_E_ GNDPWR H2 H1 H0 Net-_U63-I7_ Net-_U63-I6_ Net-_U63-I5_ VCC 74151
XU85 VCC FJ Net-_U83-Za_ Net-_U83-Zb_ Net-_U83-Zc_ Net-_U83-Zd_ VCC GNDPWR _M1VL0 FN M1V3 M1V2 M1V1 M1V0 VCC VCC NC-U85-0 NC-U85-1 NC-U85-2 74161
XU64 EPROM_2716
XU111 FS SP.A GNDPWR Net-_U111-Za_ SP.B GNDPWR Net-_U111-Zb_ GNDPWR Net-_U111-Zc_ VCC SP.C Net-_U103-D0_ VCC SP.D VCC VCC NC-U111-0 NC-U111-1 NC-U111-2 NC-U111-3 NC-U111-4 NC-U111-5 NC-U111-6 74157
XU118 VCC 7MHz GNDPWR Net-_U111-Za_ Net-_U111-Zb_ Net-_U111-Zc_ VCC GNDPWR _MHL0 VCC MH3 MH2 MH1 MH0 VCC VCC NC-U118-0 NC-U118-1 NC-U118-2 74161
XU76 VCC FJ GNDPWR GNDPWR GNDPWR GNDPWR VCC GNDPWR _M1VL0 Net-_U76-CET_ M1V7 M1V6 M1V5 M1V4 VCC VCC NC-U76-0 NC-U76-1 NC-U76-2 74161
XU91 VCC FJ Net-_U84-Za_ Net-_U84-Zb_ Net-_U84-Zc_ Net-_U84-Zd_ VCC GNDPWR _M2VL0 FN M2V3 M2V2 M2V1 M2V0 VCC VCC NC-U91-0 NC-U91-1 NC-U91-2 74161
C26 Net-_U103-TC_ GNDPWR 470p
XU103 VCC 7MHz Net-_U103-D0_ VCC GNDPWR GNDPWR VCC GNDPWR _MHL0 Net-_U103-CET_ MH7 MH6 MH5 MH4 VCC VCC NC-U103-0 NC-U103-1 NC-U103-2 74161
XU77 VCC FJ GNDPWR GNDPWR GNDPWR GNDPWR VCC GNDPWR _M2VL0 Net-_U77-CET_ M2V7 M2V6 M2V5 M2V4 VCC VCC NC-U77-0 NC-U77-1 NC-U77-2 74161
C10 _M2VL0 GNDPWR 470p
.end
