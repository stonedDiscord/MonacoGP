.title KiCad schematic
.model __D1 D
.model __D2 D
R7 Net-_IC38A-A_ VCC 100k
C19 Net-_IC38A-RCext_ Net-_IC38A-Cext_ 470m
C11 Net-_IC32B-_S_ GNDPWR 0.1m
C8 Net-_IC32B-_R_ GNDPWR 0.1m
IC32 __IC32
D1 unconnected-_D1-A-Pad2_ Net-_AE1-A_ __D1
C12 Net-_IC38A-A_ GNDPWR 0.01m
C14 Net-_IC38A-A_ GNDPWR 47
SW4 __SW4
R9 VCC Net-_IC38A-RCext_ 47k
IC33 __IC33
AE1 __AE1
RA1 __RA1
IC125 __IC125
IC37 __IC37
C3 Net-_AE1-A_ GNDPWR TILT SW.
IC12 __IC12
IC38 __IC38
IC31 __IC31
R6 VCC S-100-O 1k
R13 VCC Net-_IC49A-RCext_ 47k
C24 Net-_IC49A-RCext_ Net-_IC49A-Cext_ 100m
IC29 __IC29
IC85 __IC85
IC49 __IC49
L1 VCC Net-_TR1-C_ COIN METER
IC55 __IC55
C27 Net-_C27-Pad1_ GNDPWR 1000p
R14 Net-_IC44-Pad8_ Net-_C27-Pad1_ 220
IC44 __IC44
IC61 __IC61
R1 Net-_IC44-Pad6_ Net-_TR1-B_ 560
IC73 __IC73
TR1 __TR1
IC72 __IC72
RV1 __RV1
R5 Net-_R5-Pad1_ Net-_IC26-DIS_ R_US
IC26 __IC26
C4 Net-_IC26-CV_ GNDPWR 0.1u
D2 VCC Net-_D2-K_ __D2
R3 Net-_D2-K_ Net-_IC12-Pad8_ 220
R4 Net-_IC26-DIS_ Net-_IC26-THR_ R_US
C5 Net-_IC26-THR_ GNDPWR 77u
IC22 __IC22
C10 unconnected-_C10-Pad1_ GNDPWR 0.1m
SW2 __SW2
C7 Net-_IC32C-_R_ GNDPWR 0.1m
C6 unconnected-_C6-Pad1_ GNDPWR 0.1m
SW3 __SW3
RA2 __RA2
C9 unconnected-_C9-Pad1_ GNDPWR 0.1m
R22 VCC Net-_SW1-A_ 1k
SW1 __SW1
IC21 __IC21
IC20 __IC20
IC50 __IC50
IC74 __IC74
IC11 __IC11
IC27 __IC27
IC4 __IC4
IC16 __IC16
IC8 __IC8
IC13 __IC13
IC28 __IC28
IC10 __IC10
IC67 __IC67
IC5 __IC5
IC24 __IC24
IC17 __IC17
IC19 __IC19
IC18 __IC18
IC25 __IC25
IC79 __IC79
C41 S-100-O GNDPWR 470p
C15 Net-_IC38B-RCext_ Net-_IC38B-Cext_ 0.1m
R15 Net-_IC73-Pad12_ Net-_C25-Pad1_ 220
R8 VCC Net-_IC38B-RCext_ 47k
C25 Net-_C25-Pad1_ GNDPWR 1000p
.end
