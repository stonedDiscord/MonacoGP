.title KiCad schematic
.include "/home/stoned/MonacoGP/7400.LIB"
.include "/home/stoned/MonacoGP/IC.LIB"
.model __D2 D
.model __RV1 potentiometer( r= )
.model __D1 D
U90 __U90
U96 __U96
U97 __U97
U110 __U110
R6 VCC A30 1k
Cp36 GNDPWR VCC 100n
Cp30 GNDPWR VCC 100n
Cp32 GNDPWR VCC 100n
Cp31 GNDPWR VCC 100n
Cp38 GNDPWR VCC 100n
Cp7 GNDPWR VCC 100n
Cp9 GNDPWR VCC 100n
Cp3 GNDPWR VCC 100n
Cp5 GNDPWR VCC 100n
Cp8 GNDPWR VCC 100n
Cp21 GNDPWR VCC 100n
Cp24 GNDPWR VCC 100n
Cp27 GNDPWR VCC 100n
Cp13 GNDPWR VCC 100n
Cp29 GNDPWR VCC 100n
Cp28 GNDPWR VCC 100n
Cp26 GNDPWR VCC 100n
Cp11 GNDPWR VCC 100n
Cp4 GNDPWR VCC 100n
Cp6 GNDPWR VCC 100n
Cp12 GNDPWR VCC 100n
Cp1 GNDPWR VCC 100n
Cp19 GNDPWR VCC 100n
Cp22 GNDPWR VCC 100n
Cp14 GNDPWR VCC 100n
Cp10 GNDPWR VCC 100n
U89 __U89
Cp15 GNDPWR VCC 100n
Cp17 GNDPWR VCC 100n
Cp35 GNDPWR VCC 100n
Cp2 GNDPWR VCC 100n
Cp40 GNDPWR VCC 100n
Cp37 GNDPWR VCC 100n
Cp20 GNDPWR VCC 100n
Cp34 GNDPWR VCC 100n
Cp25 GNDPWR VCC 100n
Cp39 GNDPWR VCC 100n
Cp18 GNDPWR VCC 100n
Cp33 GNDPWR VCC 100n
Cp16 GNDPWR VCC 100n
Cp23 GNDPWR VCC 100n
U37 __U37
XU33 Net-_U33A-_R_ EXTEND__A_ Net-_U27B-Q_ VCC EXPLO.ST._G_ _EXPLO.ST._G_ 7474
U125 __U125
XU31 Net-_U20-CLR_ A26 7417
U71 __U71
U70 __U70
U95 __U95
XU73 Net-_U20-_LOAD_ Net-_U79A-MR_ 7404
U103 __U103
U104 __U104
SW1 __SW1
R22 VCC Net-_SW1-A_ 1k
XU38 Net-_U38A-A_ VCC VCC _INI._RESET__B_ unconnected-_U38B-Q-Pad5_ Net-_U38B-Cext_ Net-_U38B-RCext_ Net-_U37A-_R_ Net-_U37A-_R_ 74123
XU55 Net-_C25-Pad1_ Net-_U55-Pad11_ _EX.SIG???.??__M_ 7432
C25 Net-_C25-Pad1_ GNDPWR 1000p
R15 Net-_R15-Pad1_ Net-_C25-Pad1_ 220
R8 VCC Net-_U38B-RCext_ 47k
C15 Net-_U38B-RCext_ Net-_U38B-Cext_ 0.1m
U79 __U79
C41 A30 GNDPWR 470p
XU61 Net-_U61-Pad1_ Net-_U43B-Q_ Net-_U43A-Q_ 7402
U74 __U74
XU50 Net-_U50A-_R_ VCC _EX.SIG???.??__M_ unconnected-_U50A-_S-Pad4_ Net-_U50A-Q_ Net-_U50A-_Q_ 7474
XU22 Net-_U22-Pad1_ unconnected-_U22-Pad2_ Net-_U7-B3_ 7408
C27 Net-_C27-Pad1_ GNDPWR 1000p
C24 Net-_U49A-RCext_ Net-_U49A-Cext_ 100m
XU49 _EX.SIG???.??__M_ VCC VCC _FX.SIGNAL__B_ _SPLAY_B Net-_U49B-Cext_ Net-_U49B-RCext_ _POOL _POOL 74123
R13 VCC Net-_U49A-RCext_ 47k
XU44 Net-_U27A-Q_ Net-_U9-S1_ 7404
R14 Net-_R14-Pad1_ Net-_C27-Pad1_ 220
L1 VCC A9 COIN METER
R1 Net-_R1-Pad1_ Net-_TR1-B_ 560
TR1 __TR1
J1 __J1
U116 __U116
J3 __J3
J2 __J2
U124 __U124
U109 __U109
U117 __U117
U102 __U102
U108 __U108
U101 __U101
U75 __U75
U111 __U111
U118 __U118
XU29 Net-_U2-Pad3_ A20 7417
U57 __U57
U46 __U46
U51 __U51
C22 _LIGHT GNDPWR 470p
U56 __U56
U52 __U52
U34 __U34
U63 __U63
U119 __U119
U45 __U45
C39 Net-_U51C-_R_ GNDPWR 470p
U62 __U62
U47 __U47
U54 __U54
U80 __U80
U30 __U30
U66 __U66
SW2 __SW2
XU32 unconnected-_U32A-_R-Pad1_ Net-_U32A-_S1_ Net-_U32A-_S1_ Net-_U32A-Q_ unconnected-_U32B-_R-Pad5_ unconnected-_U32B-_S-Pad6_ Net-_U32B-Q_ 74279
R998 Net-_D2-K_ A6 220
D2 VCC Net-_D2-K_ __D2
SW3 __SW3
SW4 __SW4
XU12 Net-_U69-Za_ Net-_U10-Oa_b_ Net-_U25-UP_ 7400
ARV1 Net-_R5-Pad1_ VCC unconnected-_RV1-Pad3_ __RV1
R5 Net-_R5-Pad1_ Net-_U26-DIS_ 3.3k
C4 Net-_U26-CV_ GNDPWR 0.1u
XU26 GNDPWR Net-_U26-THR_ Net-_U26-Q_ Net-_U26-R_ Net-_U26-CV_ Net-_U26-THR_ Net-_U26-DIS_ UA555
R4 Net-_U26-DIS_ Net-_U26-THR_ 12k
C5 Net-_U26-THR_ GNDPWR 47u
U72 __U72
U21 __U21
D1 unconnected-_D1-A-Pad2_ Net-_AE1-A_ __D1
SW5 __SW5
AE1 __AE1
RA2 VCC unconnected-_RA2-R1-Pad2_ 100
R9 VCC Net-_U38A-RCext_ 47k
C19 Net-_U38A-RCext_ Net-_U38A-Cext_ 470m
C14 Net-_U38A-A_ GNDPWR 47
R7 Net-_U38A-A_ VCC 100k
C12 Net-_U38A-A_ GNDPWR 0.01m
U20 __U20
U8 __U8
U16 __U16
U27 __U27
U14 __U14
U28 __U28
U60 __U60
U18 __U18
U19 __U19
U3 __U3
C17 Net-_U40A-MR_ GNDPWR 470p
C3 Net-_U19A-MR_ GNDPWR 470p
U17 __U17
C21 Net-_U49B-RCext_ Net-_U49B-Cext_ 22m
R12 VCC Net-_U49B-RCext_ 47k
R3 VCC Net-_U1A-RCext_ 47k
U2 __U2
U40 __U40
U42 __U42
U41 __U41
U35 __U35
U36 __U36
U9 __U9
XU1 Net-_U1A-A_ Net-_U1A-B_ Net-_U1A-Clr_ Net-_U1A-_Q_ Net-_U1B-Q_ Net-_U1B-Cext_ Net-_U1B-RCext_ Net-_U1A-A_ Net-_U1A-A_ 74123
C1 Net-_U1B-RCext_ Net-_U1B-Cext_ 4.7m
C2 Net-_U1A-RCext_ Net-_U1A-Cext_ 4.7m
R2 VCC Net-_U1B-RCext_ 47k
U77 __U77
U39 __U39
U6 __U6
U4 __U4
U68 __U68
U25 __U25
U15 __U15
U69 __U69
U10 __U10
U23 __U23
U98 __U98
U76 __U76
U83 __U83
U84 __U84
U91 __U91
C26 Net-_U58-Oa=b_ GNDPWR 470p
U58 __U58
U53 __U53
U64 __U64
U65 __U65
U48 __U48
U59 __U59
C30 Net-_U119B-RCext_ Net-_U119B-Cext_ 10m
C6 PL-V-ST GNDPWR 680p
C33 Net-_U119A-RCext_ Net-_U119A-Cext_ 10m
R19 VCC Net-_U119A-RCext_ 47k
R16 VCC Net-_U119B-RCext_ 47k
U11 __U11
U24 __U24
U7 __U7
U67 __U67
U5 __U5
U13 __U13
C7 Net-_U32D-_S_ GNDPWR 0.1u
C10 unconnected-_C10-Pad1_ GNDPWR 0.1u
R10 VCC Net-_U43B-RCext_ 47k
C18 Net-_U43B-Cext_ Net-_U43B-RCext_ 15u
R11 VCC Net-_U43A-RCext_ 47k
C20 Net-_U43A-RCext_ Net-_U43A-Cext_ 10u
U43 __U43
C31 unconnected-_C31-Pad1_ unconnected-_C31-Pad2_ 100m
C32 unconnected-_C32-Pad1_ unconnected-_C32-Pad2_ 100m
XU85 Vs/16 Net-_U49A-Q_ unconnected-_U85-Pad3_ unconnected-_U85-Pad4_ 7411
.end
