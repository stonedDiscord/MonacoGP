.title KICAD
.model __RV1 potentiometer( r= )
.model __TR1 NPN level=4
.model __D1 D
J3 __J3
J2 __J2
XU73 Net-_U20-_LOAD_ Net-_U79A-MR_ 7404
XU95 Net-_U97-I6_ Net-_U85-Pad8_ Net-_U81A-_R_ 7432
XU70 Net-_U70-I3_ Net-_U70-I2_ Net-_U70-I1_ Net-_U70-I0_ unconnected-_U70-Z-Pad5_ B10 Net-_U70-_E_ GNDPWR Net-_U52B-Q2_ Net-_U52B-Q1_ Net-_U52B-Q0_ Net-_U70-I7_ Net-_U70-I6_ Net-_U70-I5_ VCC VCC NC-U70-0 NC-U70-1 NC-U70-2 74151A
XU45 Net-_U45-Pad1_ Net-_U54B-Q0_ Net-_U39B-Q1_ Net-_U39B-Q2_ 7410
XU83 7442
XU76 74153
XU61 Net-_U61-Pad1_ Net-_U43B-Q_ Net-_U43A-Q_ 7402
XU44 Net-_U27A-Q_ Net-_U9-S1_ 7404
XU68 _EXPLO._ST. BV Net-_U119A-B_ 7400
XU62 8000 BJ Net-_U62-Pad3_ 7432
XU51 Net-_U51A-_R_ Net-_U51A-_S1_ Net-_U51A-_S1_ Net-_U51A-Q_ _HOME_POS.__G_ Net-_U119A-Q_ _ACCI._ST 74279
XU48 Net-_U54B-Q2_ Net-_U54B-Q0_ Net-_U51A-_R_ 7400
XU46 Net-_U46-Pad1_ Net-_U23-Pad9_ 7404
XU77 ROM
XU47 Net-_U35-QD_ Net-_U35-QC_ NC-U47-0 Net-_U35-QB_ Net-_U35-QA_ 7420
XU36 74193
XU35 74193
XU30 Net-_U9-Zb_ Net-_U23-Pad9_ Net-_U36-DOWN_ 7400
XU91 ROM
XU84 ROM
XU65 ROM
XU56 Net-_U56-Pad1_ Net-_U64-Z_ B4 7400
XU64 Net-_U64-I3_ Net-_U64-I2_ Net-_U64-I1_ Net-_U64-I0_ Net-_U64-Z_ C15 Net-_U64-_E_ GNDPWR Net-_U52B-Q2_ Net-_U52B-Q1_ Net-_U52B-Q0_ Net-_U64-I7_ Net-_U64-I6_ Net-_U64-I5_ VCC VCC NC-U64-0 NC-U64-1 NC-U64-2 74151A
XU74 7427
C22 BC GNDPWR 470p
XU66 _ACCI. Net-_U119B-_Q_ Net-_U51C-_S1_ 7408
C26 Net-_U58-Oa=b_ GNDPWR 470p
XU58 7485
XU98 ROM
XU63 Net-_U52B-CP_ Net-_U34-Pad11_ 7MHz 7402
C39 Net-_U51C-_R_ GNDPWR 470p
XU71 ROM
XU59 ROM
XU34 Net-_U34-Pad1_ _ACCI._PULSE Net-_U27B-_S_ 7408
XU14 ACCE._C ACCE._A NC-U14-0 ACCE._B Net-_U10-B2_ 7420
XU54 74393
XU119 _SLIDE Net-_U119A-B_ VCC _SCORE_ST. SP._DOWN Net-_U119B-Cext_ Net-_U119B-RCext_ Net-_U119B-A_ Net-_U119B-A_ 74123
R16 VCC Net-_U119B-RCext_ 47k
XU72 _SP._DOWN SP._DOWN Net-_U39B-Q3_ 7402
XU39 74393
C38 B20 GNDPWR 680p
C30 Net-_U119B-RCext_ Net-_U119B-Cext_ 10m
C40 PL-V-ST. GNDPWR 680p
XU80 Net-_U10-B2_ Net-_U62-Pad3_ _ACCI._ST Net-_U14-Pad8_ 7410
XU53 7485
XU57 BD Net-_U46-Pad6_ NC-U57-0 Net-_U52A-Q1_ Net-_U52A-Q2_ 7420
C46 Net-_U59-A7_ GNDPWR 470p
C33 Net-_U119A-RCext_ Net-_U119A-Cext_ 10m
R19 VCC Net-_U119A-RCext_ 47k
C23 PL-H-ST. GNDPWR 470p
XU52 74393
XU97 Net-_U100A-1Y_ Net-_U90-Q0_ Net-_RA3-R4_ Net-_U90-Q1_ Net-_RA3-R3_ Net-_U90-Q2_ Net-_RA3-R2_ GNDPWR Net-_RA3-R1_ Net-_U90-Q3_ unconnected-_U97-O5b-Pad11_ unconnected-_U97-I5-Pad12_ Net-_RA3-R5_ Net-_U97-I6_ VCC VCC NC-U97-0 NC-U97-1 NC-U97-2 NC-U97-3 74367A
XU100 Net-_U100A-1A_ Net-_U100B-2A_ AREA_5 Net-_U100B-2C_ AREA_2 Net-_U100B-2Y_ GNDPWR Net-_U100A-1Y_ Net-_U100A-1C_ AREA_4 unconnected-_U100A-1X-Pad11_ unconnected-_U100A-1_X-Pad12_ VCC VCC NC-U100-0 NC-U100-1 NC-U100-2 7450
XU110 Net-_U100B-2Y_ Net-_U104-Q0_ Net-_RA3-R4_ Net-_U104-Q1_ Net-_RA3-R3_ Net-_U104-Q2_ Net-_RA3-R2_ GNDPWR Net-_RA3-R1_ Net-_U104-Q3_ unconnected-_U110-O5b-Pad11_ unconnected-_U110-I5-Pad12_ Net-_RA3-R5_ Net-_U110-I6_ VCC VCC NC-U110-0 NC-U110-1 NC-U110-2 NC-U110-3 74367A
XU122 Net-_U122-Pad1_ Net-_U109-Q2_ Net-_U109-Q0_ 7402
XU123 Net-_U96-Q1_ Net-_U96-Q3_ Net-_U109-Q1_ Net-_U122-Pad1_ 7410
XU90 VCC Net-_U101-_PE_ Net-_U89-Za_ Net-_U89-Zb_ Net-_U89-Zc_ Net-_U89-Zd_ VCC GNDPWR Net-_U90-_PE_ CN Net-_U90-Q3_ Net-_U90-Q2_ Net-_U90-Q1_ Net-_U90-Q0_ VCC VCC NC-U90-0 NC-U90-1 NC-U90-2 74161
XU82 Net-_U117-D3_ Net-_U117-D1_ 7404
XU96 VCC Net-_U101-_PE_ GNDPWR GNDPWR GNDPWR GNDPWR VCC GNDPWR Net-_U90-_PE_ Net-_U90-TC_ Net-_U96-Q3_ Net-_U96-Q2_ Net-_U96-Q1_ Net-_U96-Q0_ VCC VCC NC-U96-0 NC-U96-1 NC-U96-2 74161
XU89 Net-_U89-S_ GNDPWR VCC Net-_U89-Za_ GNDPWR Net-_U89-I1b_ Net-_U89-Zb_ GNDPWR Net-_U89-Zc_ Net-_U89-I1b_ GNDPWR Net-_U89-Zd_ Net-_U121A-B_ VCC VCC VCC NC-U89-0 NC-U89-1 NC-U89-2 NC-U89-3 NC-U89-4 NC-U89-5 NC-U89-6 74157
XU99 VCC Net-_U105-D1_ Net-_U99A-C_ VCC Net-_U100A-1A_ unconnected-_U99A-_Q-Pad6_ 7474
XU93 Net-_U100A-1B_ Net-_U66-Pad4_ Net-_U99A-C_ 7408
XU86 unconnected-_U86-Pad1_ unconnected-_U86-Pad2_ unconnected-_U86-Pad3_ 7402
XU107 Net-_U121A-Q_ Net-_U107-Pad2_ Net-_U87B-Q_ Net-_U101-Q1_ 7410
XU104 VCC Net-_U101-_PE_ Net-_U103-Za_ Net-_U103-Zb_ Net-_U103-Zc_ Net-_U103-Zd_ VCC GNDPWR Net-_U104-_PE_ CN Net-_U104-Q3_ Net-_U104-Q2_ Net-_U104-Q1_ Net-_U104-Q0_ VCC VCC NC-U104-0 NC-U104-1 NC-U104-2 74161
XU103 Net-_U103-S_ GNDPWR VCC Net-_U103-Za_ GNDPWR Net-_U103-I1b_ Net-_U103-Zb_ GNDPWR Net-_U103-Zc_ Net-_U103-I1b_ GNDPWR Net-_U103-Zd_ Net-_U103-I1d_ VCC VCC VCC NC-U103-0 NC-U103-1 NC-U103-2 NC-U103-3 NC-U103-4 NC-U103-5 NC-U103-6 74157
XU117 VCC Net-_U101-_PE_ VCC Net-_U117-D1_ Net-_U117-D1_ Net-_U117-D3_ VCC GNDPWR Net-_U116-_PE_ CN Net-_U117-Q3_ Net-_U117-Q2_ Net-_U117-Q1_ Net-_U117-Q0_ VCC VCC NC-U117-0 NC-U117-1 NC-U117-2 74161
XU109 VCC Net-_U101-_PE_ GNDPWR GNDPWR GNDPWR GNDPWR VCC GNDPWR Net-_U104-_PE_ Net-_U104-TC_ Net-_U109-Q3_ Net-_U109-Q2_ Net-_U109-Q1_ Net-_U109-Q0_ VCC VCC NC-U109-0 NC-U109-1 NC-U109-2 74161
XU114 Net-_U118-Zb_ BS 7404
XU81 Net-_U81A-_R_ Net-_U81A-_S1_ Net-_U81A-_S1_ Net-_U121A-B_ Net-_U81B-_R_ Net-_U81B-_S_ Net-_U117-D3_ 74279
XU105 74S288
XU92 VCC Net-_U105-D2_ Net-_U92A-C_ VCC Net-_U100B-2C_ unconnected-_U92A-_Q-Pad6_ 7474
C29 Net-_U112A-CP_ GNDPWR 470m
XU124 Net-_U124-OEa_ Net-_U117-Q0_ Net-_RA3-R4_ Net-_U117-Q1_ Net-_RA3-R3_ Net-_U117-Q2_ Net-_RA3-R2_ GNDPWR Net-_RA3-R1_ Net-_U117-Q3_ unconnected-_U124-O5b-Pad11_ unconnected-_U124-I5-Pad12_ Net-_RA3-R5_ Net-_U124-I6_ VCC VCC NC-U124-0 NC-U124-1 NC-U124-2 NC-U124-3 74367A
XU21 74192
XU20 74192
XU125 unconnected-_U125-Pad1_ unconnected-_U125-Pad2_ Net-_SW1-B_ Net-_U32A-Q_ 7411
XU32 Net-_U32A-_R_ Net-_RN2C-R3.1_ Net-_RN2C-R3.1_ Net-_U32A-Q_ Net-_RN2D-R4.1_ Net-_RN2E-R5.1_ Net-_U32B-Q_ 74279
RN2 Net-_RN2A-R1.1_ Net-_RN2B-R2.1_ 100
C36 Net-_RN2G-R7.2_ GNDPWR 0.1m
XU37 Net-_U37A-_R_ VCC Net-_U20-_LOAD_ VCC B1 BD 7474
XU33 Net-_U33A-_R_ BB Net-_U27B-Q_ unconnected-_U33A-_S-Pad4_ EXPLO._ST. _EXPLO._ST. 7474
XU12 Net-_U69-Za_ Net-_U10-Oa_b_ Net-_U25-UP_ 7400
XU22 Net-_U22-Pad1_ Net-_U32D-Q_ Net-_U7-B3_ 7408
XU26 GNDPWR Net-_U26-THR_ Net-_U26-Q_ Net-_U26-R_ Net-_U26-CV_ Net-_U26-THR_ Net-_U26-DIS_ UA555
C4 Net-_U26-CV_ GNDPWR 0.1u
C5 Net-_U26-THR_ GNDPWR 47u
R5 Net-_R5-Pad1_ Net-_U26-DIS_ 3.3k
R4 Net-_U26-DIS_ Net-_U26-THR_ 12k
ARV1 Net-_R5-Pad1_ VCC unconnected-_RV1-Pad3_ __RV1
XU31 Net-_U20-CLR_ A26 7417
R24 A32 Net-_U32C-_R_ 100
R23 VCC A32 560
R6 VCC A30 1k
R1 Net-_R1-Pad1_ Net-_TR1-B_ 560
QTR1 Net-_TR1-B_ A9 GNDPWR __TR1
C37 Net-_U32C-_R_ GNDPWR 0.1m
C8 Net-_RN2C-R3.1_ GNDPWR 0.1u
C11 Net-_U32A-_R_ GNDPWR 470m
C9 Net-_RN2E-R5.1_ GNDPWR 0.1u
SW1 __SW1
R22 VCC Net-_SW1-A_ 1k
C12 Net-_RN2H-R8.1_ GNDPWR 0.01m
R7 Net-_RN2H-R8.1_ VCC 100k
D1 Net-_D1-A_ Aj __D1
C6 Net-_RN2D-R4.1_ GNDPWR 680p
R9 VCC Net-_U38A-RCext_ 47k
C19 Net-_U38A-RCext_ Net-_U38A-Cext_ 470m
XU38 Net-_RN2H-R8.1_ VCC VCC Ak unconnected-_U38B-Q-Pad5_ Net-_U38B-Cext_ Net-_U38B-RCext_ Net-_U37A-_R_ Net-_U37A-_R_ 74123
C13 Net-_RN2H-R8.1_ Net-_RN2H-R8.1_ 0.01m
C14 Net-_RN2H-R8.1_ GNDPWR 47
C32 Net-_U121B-RCext_ Net-_U121B-Cext_ 470m
R18 VCC Net-_U121B-RCext_ 47k
C34 Net-_U120A-RCext_ Net-_U120A-Cext_ 470m
R20 Net-_U120A-RCext_ VCC 47k
XU121 Net-_U121A-A_ Net-_U121A-B_ BRIDGE_AP. Net-_U121A-_Q_ Net-_U121A-A_ Net-_U121B-Cext_ Net-_U121B-RCext_ Net-_U121A-B_ Net-_U121A-B_ 74123
XU88 Net-_U85-Pad6_ Net-_U110-I6_ Net-_U81D-_S_ 7432
XU85 B21 Net-_U49A-Q_ unconnected-_U85-Pad3_ CC 7411
R21 VCC Net-_U121A-RCext_ 47k
C35 Net-_U121A-RCext_ Net-_U121A-Cext_ 470m
Cp17 GNDPWR VCC 100n
Cp29 GNDPWR VCC 100n
Cp12 GNDPWR VCC 100n
Cp30 GNDPWR VCC 100n
Cp22 GNDPWR VCC 100n
Cp34 GNDPWR VCC 100n
Cp23 GNDPWR VCC 100n
Cp9 GNDPWR VCC 100n
Cp5 GNDPWR VCC 100n
Cp2 GNDPWR VCC 100n
Cp8 GNDPWR VCC 100n
Cp3 GNDPWR VCC 100n
Cp1 GNDPWR VCC 100n
Cp4 GNDPWR VCC 100n
Cp46 GNDPWR VCC 100n
Cp27 GNDPWR VCC 100n
Cp32 GNDPWR VCC 100n
Cp14 GNDPWR VCC 100n
Cp31 GNDPWR VCC 100n
Cp42 GNDPWR VCC 100n
Cp20 GNDPWR VCC 100n
Cp33 GNDPWR VCC 100n
Cp13 GNDPWR VCC 100n
Cp7 GNDPWR VCC 100n
Cp6 GNDPWR VCC 100n
Cp16 GNDPWR VCC 100n
Cp41 GNDPWR VCC 100n
Cp18 GNDPWR VCC 100n
Cp11 GNDPWR VCC 100n
Cp15 GNDPWR VCC 100n
Cp26 GNDPWR VCC 100n
Cp43 GNDPWR VCC 100n
Cp28 GNDPWR VCC 100n
Cp37 GNDPWR VCC 100n
Cp40 GNDPWR VCC 100n
Cp36 GNDPWR VCC 100n
Cp35 GNDPWR VCC 100n
Cp38 GNDPWR VCC 100n
Cp10 GNDPWR VCC 100n
Cp19 GNDPWR VCC 100n
Cp39 GNDPWR VCC 100n
Cp25 GNDPWR VCC 100n
Cp47 GNDPWR VCC 100n
Cp24 GNDPWR VCC 100n
Cp21 GNDPWR VCC 100n
Cp44 GNDPWR VCC 100n
Cp45 GNDPWR VCC 100n
Cp48 GNDPWR VCC 100n
XU49 B2 VCC VCC C1 _SPLAY_B Net-_U49B-Cext_ Net-_U49B-RCext_ CM CM 74123
C24 Net-_U49A-RCext_ Net-_U49A-Cext_ 100m
XU55 Net-_C25-Pad1_ Net-_U55-Pad11_ B2 7432
XU50 Net-_U50A-_R_ VCC B2 unconnected-_U50A-_S-Pad4_ Net-_U50A-Q_ Net-_U50A-_Q_ 7474
C27 Net-_C27-Pad1_ GNDPWR 1000p
R14 Net-_R14-Pad1_ Net-_C27-Pad1_ 220
R13 VCC Net-_U49A-RCext_ 47k
R15 Net-_R15-Pad1_ Net-_C25-Pad1_ 220
C25 Net-_C25-Pad1_ GNDPWR 1000p
C143 A30 GNDPWR 470p
XU79 74393
R8 VCC Net-_U38B-RCext_ 47k
C15 Net-_U38B-RCext_ Net-_U38B-Cext_ 0.1m
C66 Net-_U75A-C_ GNDPWR 470m
XU106 Net-_U106-Pad1_ Net-_U101-Q3_ AREA_4 7408
XU112 74393
C43 Net-_U124-OEa_ GNDPWR 470m
XU75 VCC Net-_U75A-D_ Net-_U75A-C_ VCC Net-_U75A-Q_ unconnected-_U75A-_Q-Pad6_ 7474
C28 Net-_U100A-1B_ GNDPWR 470m
XU94 Net-_U101-Q1_ Net-_U101-Q2_ Net-_U101-Q3_ AREA_2 unconnected-_U94-Q1-Pad5_ unconnected-_U94-Q2-Pad6_ unconnected-_U94-Q3-Pad7_ GNDPWR Net-_U100A-1B_ AREA_1 unconnected-_U94-Q6-Pad11_ AREA_5 VCC Net-_U87B-_Q_ VCC VCC NC-U94-0 NC-U94-1 NC-U94-2 NC-U94-3 NC-U94-4 NC-U94-5 74259
XU102 VCC 7MHz Net-_U102-D0_ Net-_U102-D1_ Net-_U102-D2_ Net-_U102-D3_ Net-_U102-CEP_ GNDPWR Net-_U101-_PE_ VCC Net-_U102-Q3_ Net-_U102-Q2_ Net-_U102-Q1_ Net-_U102-Q0_ VCC VCC NC-U102-0 NC-U102-1 NC-U102-2 74161
XU116 VCC Net-_U101-_PE_ GNDPWR GNDPWR GNDPWR GNDPWR VCC GNDPWR Net-_U116-_PE_ Net-_U116-CET_ Net-_U116-Q3_ Net-_U116-Q2_ Net-_U116-Q1_ Net-_U116-Q0_ VCC VCC NC-U116-0 NC-U116-1 NC-U116-2 74161
C42 Net-_U101-TC_ GNDPWR 470p
XU87 unconnected-_U87A-J-Pad1_ unconnected-_U87A-_Q-Pad2_ unconnected-_U87A-Q-Pad3_ unconnected-_U87A-K-Pad4_ Net-_U87B-Q_ Net-_U87B-_Q_ VCC VCC 74107
XU101 VCC 7MHz VCC VCC GNDPWR GNDPWR VCC GNDPWR Net-_U101-_PE_ Net-_U101-CET_ Net-_U101-Q3_ Net-_U101-Q2_ Net-_U101-Q1_ Net-_U101-Q0_ VCC VCC NC-U101-0 NC-U101-1 NC-U101-2 74161
XU118 Net-_U102-Q0_ Net-_U111-D0_ Net-_U111-D1_ unconnected-_U118-Za-Pad4_ Net-_U111-D2_ Net-_U111-D3_ Net-_U118-Zb_ GNDPWR Net-_U118-Zc_ Net-_U111-D5_ Net-_U111-D4_ Net-_U118-Zd_ Net-_U111-D7_ Net-_U111-D6_ VCC VCC NC-U118-0 NC-U118-1 NC-U118-2 NC-U118-3 NC-U118-4 NC-U118-5 NC-U118-6 74157
C45 Net-_U118-Zb_ GNDPWR 470p
XU111 ROM
XU29 Net-_U2-Pad3_ A20 7417
XU120 Net-_U120A-A_ Net-_U103-I1d_ BRIDGE_AP. Net-_U120A-_Q_ Net-_U120A-A_ Net-_U120B-Cext_ Net-_U120B-RCext_ Net-_U103-I1d_ Net-_U103-I1d_ 74123
C31 Net-_U120B-RCext_ Net-_U120B-Cext_ 470m
R17 VCC Net-_U120B-RCext_ 47k
XU40 74393
V1 VCC GNDPWR DC 1 
XU113 7485
C86 Ah GNDPWR 0.01m
XU115 74S288
XU108 CS Net-_U108-I0a_ GNDPWR Net-_U102-D0_ Net-_U108-I0b_ GNDPWR Net-_U102-D1_ GNDPWR Net-_U102-D2_ GNDPWR Net-_U108-I0c_ Net-_U102-D3_ VCC Net-_U108-I0d_ VCC VCC NC-U108-0 NC-U108-1 NC-U108-2 NC-U108-3 NC-U108-4 NC-U108-5 NC-U108-6 74157
R11 VCC Net-_U43A-RCext_ 47k
C20 Net-_U43A-RCext_ Net-_U43A-Cext_ 10u
XU43 CA PLAYER Net-_U15-QD_ Net-_U1A-A_ Net-_U43B-Q_ Net-_U43B-Cext_ Net-_U43B-RCext_ CM CM 74123
C18 Net-_U43B-Cext_ Net-_U43B-RCext_ 15u
R10 VCC Net-_U43B-RCext_ 47k
C21 Net-_U49B-RCext_ Net-_U49B-Cext_ 22m
R12 VCC Net-_U49B-RCext_ 47k
C1 Net-_U1B-RCext_ Net-_U1B-Cext_ 4.7m
XU2 Net-_U3-S0_ _SP._DOWN Net-_U2-Pad3_ 7408
XU1 Net-_U1A-A_ A8 Net-_U1A-Clr_ Net-_U1A-_Q_ Net-_U1B-Q_ Net-_U1B-Cext_ Net-_U1B-RCext_ Net-_U1A-A_ Net-_U1A-A_ 74123
C2 Net-_U1A-RCext_ Net-_U1A-Cext_ 4.7m
R2 VCC Net-_U1B-RCext_ 47k
R3 VCC Net-_U1A-RCext_ 47k
XU60 Net-_U60-S_ B21 BX Net-_U60-Za_ B22 Vs/8 Net-_U60-Zb_ GNDPWR unconnected-_U60-Zc-Pad9_ unconnected-_U60-I1c-Pad10_ unconnected-_U60-I0c-Pad11_ unconnected-_U60-Zd-Pad12_ unconnected-_U60-I1d-Pad13_ unconnected-_U60-I0d-Pad14_ VCC VCC NC-U60-0 NC-U60-1 NC-U60-2 NC-U60-3 NC-U60-4 NC-U60-5 NC-U60-6 74157
C44 C12 GNDPWR 470p
XU78 74393
XU28 unconnected-_U28-Pad1_ unconnected-_U28-Pad2_ Net-_U10-A1_ Net-_U10-A0_ 7410
XU27 Net-_U27A-_R_ Net-_U27A-_S1_ Net-_U27A-_S1_ Net-_U27A-Q_ _HOME_POS.__G_ Net-_U27B-_S_ Net-_U27B-Q_ 74279
XU23 EXPLO._ST. Net-_U27B-Q_ Net-_U27A-_R_ 7432
XU16 VCC Net-_U27A-_R_ _ACCI. 7486
C16 Net-_U39A-CP_ GNDPWR 470p
XU13 ACCE._D A12 7407
C7 Net-_RN2A-R1.1_ GNDPWR 0.1u
XU6 Net-_U15-QD_ Net-_U10-B2_ 7404
C10 Net-_RN2B-R2.1_ GNDPWR 0.1u
XU19 74393
XU69 74153
XU24 74193
XU11 7485
XU67 B12 B12 Net-_U67B-2B_ BN Net-_U67B-2D_ Net-_U5A-CP_ GNDPWR Net-_U67A-1Y_ BN Net-_U67A-1D_ unconnected-_U67A-1X-Pad11_ unconnected-_U67A-1_X-Pad12_ VCC VCC NC-U67-0 NC-U67-1 NC-U67-2 7450
XU10 7485
XU5 74393
XU8 Vs/8 Net-_U7-Oa_b_ Net-_U15-DOWN_ 7400
XU7 7485
XU15 74193
XU4 Net-_U4-I2_ Net-_U4-I2_ Net-_U4-I0_ Net-_U4-I0_ Net-_U4-Z_ unconnected-_U4-_Z-Pad6_ Net-_U27A-_R_ GNDPWR Net-_U10-B2_ Net-_U10-B1_ Net-_U10-B0_ Net-_U4-I6_ Net-_U4-I6_ Net-_U4-I4_ VCC VCC NC-U4-0 NC-U4-1 NC-U4-2 74151A
C17 Net-_U40A-MR_ GNDPWR 470p
C3 Net-_U19A-MR_ GNDPWR 470p
XU9 74153
XU3 74153
XU18 7485
XU42 7485
XU25 74193
XU41 7485
XU17 7485
C41 Net-_U101-_PE_ GNDPWR 470p
J1 __J1
.end
