.title KiCad schematic
.model __D1 D
.model __D3 D
.model __D2 D
Cp28 GNDPWR VCC C
Cp10 GNDPWR VCC C
Cp17 GNDPWR VCC C
Cp9 GNDPWR VCC C
Cp5 GNDPWR VCC C
Cp30 GNDPWR VCC C
Cp33 GNDPWR VCC C
Cp34 GNDPWR VCC C
Cp20 GNDPWR VCC C
Cp19 GNDPWR VCC C
Cp22 GNDPWR VCC C
Cp36 GNDPWR VCC C
Cp31 GNDPWR VCC C
Cp21 GNDPWR VCC C
Cp35 GNDPWR VCC C
Cp27 GNDPWR VCC C
Cp32 GNDPWR VCC C
Cp29 GNDPWR VCC C
Cp2 GNDPWR VCC C
Cp13 GNDPWR VCC C
Cp1 GNDPWR VCC C
Cp15 GNDPWR VCC C
Cp4 GNDPWR VCC C
Cp16 GNDPWR VCC C
Cp14 GNDPWR VCC C
Cp12 GNDPWR VCC C
Cp7 GNDPWR VCC C
Cp8 GNDPWR VCC C
Cp18 GNDPWR VCC C
Cp6 GNDPWR VCC C
Cp11 GNDPWR VCC C
Cp3 GNDPWR VCC C
Cp24 GNDPWR VCC C
Cp25 GNDPWR VCC C
Cp26 GNDPWR VCC C
Cp23 GNDPWR VCC C
U31 __U31
U45 __U45
U201 __U201
U22 __U22
U9 __U9
U86 __U86
U1 __U1
U15 __U15
U4 __U4
U8 __U8
U3 __U3
U21 __U21
U19 __U19
U44 __U44
U66 __U66
U7 __U7
U13 __U13
U14 __U14
J2 __J2
U18 __U18
U23 __U23
J1 __J1
U56 __U56
U59 __U59
U50 __U50
U65 __U65
U52 __U52
U10 __U10
U12 __U12
U17 __U17
U27 __U27
U26 __U26
U34 __U34
U58 __U58
U2 __U2
U79 __U79
U20 __U20
U5 __U5
U40 __U40
C2 Net-_U40B-_Q_ GNDPWR 470p
U49 __U49
U39 __U39
U48 __U48
U41 __U41
U33 __U33
U32 __U32
U47 __U47
C1 _COIN_IN GNDPWR 470p
U25 __U25
Q1 __Q1
R13 GNDPWR D11 10k
R1 VCC D11 470
R6 Net-_R6-Pad1_ D13 470
D1 D11 Net-_D1-K_ __D1
D3 D13 Net-_D1-K_ __D3
D2 D12 Net-_D1-K_ __D2
R5 VCC D13 470
R3 VCC D12 470
R4 Net-_R4-Pad1_ D12 470
R2 Net-_R2-Pad1_ D11 470
R14 GNDPWR D12 10k
R15 GNDPWR D13 10k
U72 __U72
U67 __U67
RN1 __RN1
U75 __U75
U82 __U82
U89 __U89
U38 __U38
U88 __U88
U43 __U43
U42 __U42
U202 __U202
U28 __U28
U37 __U37
U35 __U35
U36 __U36
U57 __U57
U62 __U62
U60 __U60
U55 __U55
U61 __U61
U29 __U29
U24 __U24
U30 __U30
U73 __U73
U46 __U46
U53 __U53
U51 __U51
U16 __U16
U11 __U11
U6 __U6
U69 __U69
U70 __U70
U84 __U84
U85 __U85
U76 __U76
U54 __U54
U83 __U83
U68 __U68
U91 __U91
U77 __U77
U63 __U63
U71 __U71
U64 __U64
U78 __U78
U90 __U90
U80 __U80
U81 __U81
U87 __U87
U74 __U74
.end
