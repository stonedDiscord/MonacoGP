.title KiCad schematic
.include "/home/stoned/MonacoGP/7400.LIB"
.include "/home/stoned/MonacoGP/IC.LIB"
.model __RV1 potentiometer( r= )
.model __D2 D
.model __D1 D
.model __TR1 NPN level=4
C39 Net-_U51C-_R_ GNDPWR 470p
XU56 Net-_U56-Pad1_ Net-_U64-Z_ B4 7400
XU51 Net-_U51A-_R_ Net-_U51A-_S1_ Net-_U51A-_S1_ Net-_U51A-Q_ _HOME_POS.__G_ Net-_U119A-Q_ _ACCI._ST 74279
C26 Net-_U58-Oa=b_ GNDPWR 470p
U58 U58.unbekannt
XU66 _ACCI. Net-_U119B-_Q_ Net-_U51C-_S1_ 7408
XU62 8000 BZ Net-_U62-Pad3_ 7432
XU57 _COIN_IN Net-_U46-Pad6_ NC-U57-0 Net-_U52A-Q1_ Net-_U52A-Q2_ 7420
U53 __U53
XU119 _SLIDE Net-_U119A-B_ VCC _SCORE_ST. SP._DOWN Net-_U119B-Cext_ Net-_U119B-RCext_ Net-_U119B-A_ Net-_U119B-A_ 74123
C33 Net-_U119A-RCext_ Net-_U119A-Cext_ 10m
R19 VCC Net-_U119A-RCext_ 47k
U59 __U59
XU46 Net-_U46-Pad1_ Net-_U23-Pad9_ 7404
J2 __J2
J1 __J1
U64 __U64
XU54 74393
XU48 Net-_U54B-Q2_ Net-_U54B-Q0_ Net-_U51A-_R_ 7400
XU72 _SP._DOWN SP._DOWN Net-_U39B-Q3_ 7402
XU45 Net-_U45-Pad1_ Net-_U54B-Q0_ Net-_U39B-Q1_ Net-_U39B-Q2_ 7410
R16 VCC Net-_U119B-RCext_ 47k
C30 Net-_U119B-RCext_ Net-_U119B-Cext_ 10m
U39 U39.unbekannt
C38 B20 GNDPWR 680p
U91 __U91
U98 __U98
XU44 Net-_U27A-Q_ Net-_U9-S1_ 7404
XU63 Net-_U52B-CP_ Net-_U34-Pad11_ 7MHz 7402
C22 _LIGHT GNDPWR 470p
U84 __U84
U65 __U65
XU74 7427
U71 __U71
XU70 Net-_U70-I3_ Net-_U70-I2_ Net-_U70-I1_ Net-_U70-I0_ unconnected-_U70-Z-Pad5_ B10 Net-_U70-_E_ GNDPWR Net-_U52B-Q2_ Net-_U52B-Q1_ Net-_U52B-Q0_ Net-_U70-I7_ Net-_U70-I6_ Net-_U70-I5_ VCC VCC NC-U70-0 NC-U70-1 NC-U70-2 74151A
J3 __J3
U83 U83.unbekannt
U76 U76.unbekannt
XU61 Net-_U61-Pad1_ Net-_U43B-Q_ Net-_U43A-Q_ 7402
XU68 _EXPLO._ST. _PLAYER_BODY Net-_U119A-B_ 7400
XU73 Net-_U20-_LOAD_ Net-_U79A-MR_ 7404
XU95 Net-_U97-I6_ Net-_U85-Pad8_ Net-_U81A-_R_ 7432
XU30 Net-_U9-Zb_ Net-_U23-Pad9_ Net-_U36-DOWN_ 7400
XU47 Net-_U35-QD_ Net-_U35-QC_ NC-U47-0 Net-_U35-QB_ Net-_U35-QA_ 7420
U52 __U52
XU34 Net-_U34-Pad1_ _ACCI._PULSE Net-_U27B-_S_ 7408
XU80 EXT.CAR_CONT. Net-_U62-Pad3_ _ACCI._ST Net-_U14-Pad8_ 7410
C40 PL-V-ST GNDPWR 680p
XU112 74393
XU123 Net-_U96-Q1_ Net-_U96-Q3_ Net-_U109-Q1_ Net-_U122-Pad1_ 7410
XU92 VCC Net-_U105-D2_ Net-_U92A-C_ VCC Net-_U100B-2C_ unconnected-_U92A-_Q-Pad6_ 7474
XU100 Net-_U100A-1A_ Net-_U100B-2A_ AREA_5 Net-_U100B-2C_ AREA_2 Net-_U100B-2Y_ GNDPWR Net-_U100A-1Y_ Net-_U100A-1C_ AREA_4 unconnected-_U100A-1X-Pad11_ unconnected-_U100A-1_X-Pad12_ VCC VCC NC-U100-0 NC-U100-1 NC-U100-2 7450
XU114 Net-_U118-Zb_ _OTHER_TIRE 7404
XU87 unconnected-_U87A-J-Pad1_ unconnected-_U87A-_Q-Pad2_ unconnected-_U87A-Q-Pad3_ unconnected-_U87A-K-Pad4_ Net-_U87B-Q_ Net-_U87B-_Q_ VCC VCC 74107
XU93 AREA_3 Net-_U66-Pad4_ Net-_U99A-C_ 7408
XU122 Net-_U122-Pad1_ Net-_U109-Q2_ Net-_U109-Q0_ 7402
XU75 VCC Net-_U75A-D_ Net-_U75A-C_ VCC Net-_U75A-Q_ unconnected-_U75A-_Q-Pad6_ 7474
XU118 Net-_U102-Q0_ Net-_U111-D0_ Net-_U111-D1_ unconnected-_U118-Za-Pad4_ Net-_U111-D2_ Net-_U111-D3_ Net-_U118-Zb_ GNDPWR Net-_U118-Zc_ Net-_U101-Q0_ Net-_U111-D4_ Net-_U118-Zd_ Net-_U101-Q0_ Net-_U111-D6_ VCC VCC NC-U118-0 NC-U118-1 NC-U118-2 NC-U118-3 NC-U118-4 NC-U118-5 NC-U118-6 74157
XU124 Net-_U124-OEa_ Net-_U117-Q0_ Net-_RA3-R4_ Net-_U117-Q1_ Net-_RA3-R3_ Net-_U117-Q2_ Net-_RA3-R2_ GNDPWR Net-_RA3-R1_ Net-_U117-Q3_ unconnected-_U124-O5b-Pad11_ unconnected-_U124-I5-Pad12_ Net-_RA3-R5_ Net-_U124-I6_ VCC VCC NC-U124-0 NC-U124-1 NC-U124-2 NC-U124-3 74367A
XU110 Net-_U100B-2Y_ Net-_U104-Q0_ Net-_RA3-R4_ Net-_U104-Q1_ Net-_RA3-R3_ Net-_U104-Q2_ Net-_RA3-R2_ GNDPWR Net-_RA3-R1_ Net-_U104-Q3_ unconnected-_U110-O5b-Pad11_ unconnected-_U110-I5-Pad12_ Net-_RA3-R5_ Net-_U110-I6_ VCC VCC NC-U110-0 NC-U110-1 NC-U110-2 NC-U110-3 74367A
XU97 Net-_U100A-1Y_ Net-_U90-Q0_ Net-_RA3-R4_ Net-_U90-Q1_ Net-_RA3-R3_ Net-_U90-Q2_ Net-_RA3-R2_ GNDPWR Net-_RA3-R1_ Net-_U90-Q3_ unconnected-_U97-O5b-Pad11_ unconnected-_U97-I5-Pad12_ Net-_RA3-R5_ Net-_U97-I6_ VCC VCC NC-U97-0 NC-U97-1 NC-U97-2 NC-U97-3 74367A
XU101 VCC 7MHz VCC VCC GNDPWR GNDPWR VCC GNDPWR Net-_U101-_PE_ Net-_U101-CET_ Net-_U101-Q3_ Net-_U101-Q2_ Net-_U101-Q1_ Net-_U101-Q0_ VCC VCC NC-U101-0 NC-U101-1 NC-U101-2 74161
U78 U78.unbekannt
XU106 Net-_U106-Pad1_ Net-_U101-Q3_ AREA_4 7408
C42 Net-_U124-OEa_ GNDPWR 470m
U111 __U111
XU108 Net-_U108-S_ Net-_U108-I0a_ GNDPWR Net-_U102-D0_ Net-_U108-I0b_ GNDPWR Net-_U102-D1_ GNDPWR Net-_U102-D2_ GNDPWR Net-_U108-I0c_ Net-_U102-D3_ VCC Net-_U108-I0d_ VCC VCC NC-U108-0 NC-U108-1 NC-U108-2 NC-U108-3 NC-U108-4 NC-U108-5 NC-U108-6 74157
XU107 Net-_U121A-Q_ Net-_U107-Pad2_ Net-_U87B-Q_ Net-_U101-Q1_ 7410
XU94 Net-_U101-Q1_ Net-_U101-Q2_ Net-_U101-Q3_ AREA_2 unconnected-_U94-Q1-Pad5_ unconnected-_U94-Q2-Pad6_ unconnected-_U94-Q3-Pad7_ GNDPWR AREA_3 AREA_1 unconnected-_U94-Q6-Pad11_ AREA_5 VCC Net-_U87B-_Q_ VCC VCC NC-U94-0 NC-U94-1 NC-U94-2 NC-U94-3 NC-U94-4 NC-U94-5 74259
C28 AREA_3 GNDPWR 470m
C29 Net-_U112A-CP_ GNDPWR 470m
XU86 unconnected-_U86-Pad1_ unconnected-_U86-Pad2_ unconnected-_U86-Pad3_ 7402
U105 __U105
C66 Net-_U75A-C_ GNDPWR 470m
XU82 Net-_U117-D3_ Net-_U117-D1_ 7404
XU99 VCC Net-_U105-D1_ Net-_U99A-C_ VCC Net-_U100A-1A_ unconnected-_U99A-_Q-Pad6_ 7474
XU96 VCC Net-_U101-_PE_ GNDPWR GNDPWR GNDPWR GNDPWR VCC GNDPWR Net-_U90-_PE_ Net-_U90-TC_ Net-_U96-Q3_ Net-_U96-Q2_ Net-_U96-Q1_ Net-_U96-Q0_ VCC VCC NC-U96-0 NC-U96-1 NC-U96-2 74161
XU104 VCC Net-_U101-_PE_ Net-_U103-Za_ Net-_U103-Zb_ Net-_U103-Zc_ Net-_U103-Zd_ VCC GNDPWR Net-_U104-_PE_ _Vb Net-_U104-Q3_ Net-_U104-Q2_ Net-_U104-Q1_ Net-_U104-Q0_ VCC VCC NC-U104-0 NC-U104-1 NC-U104-2 74161
XU103 Net-_U103-S_ GNDPWR VCC Net-_U103-Za_ GNDPWR Net-_U103-I1b_ Net-_U103-Zb_ GNDPWR Net-_U103-Zc_ Net-_U103-I1b_ GNDPWR Net-_U103-Zd_ Net-_U103-I1d_ VCC VCC VCC NC-U103-0 NC-U103-1 NC-U103-2 NC-U103-3 NC-U103-4 NC-U103-5 NC-U103-6 74157
XU88 Net-_U85-Pad6_ Net-_U110-I6_ Net-_U81D-_S_ 7432
XU81 Net-_U81A-_R_ Net-_U81A-_S1_ Net-_U81A-_S1_ Net-_U121A-B_ Net-_U81B-_R_ Net-_U81B-_S_ Net-_U117-D3_ 74279
U113 U113.unbekannt
XU120 Net-_U120A-A_ Net-_U103-I1d_ Net-_U120A-Clr_ Net-_U120A-_Q_ Net-_U120A-A_ Net-_U120B-Cext_ Net-_U120B-RCext_ Net-_U103-I1d_ Net-_U103-I1d_ 74123
R20 Net-_U120A-RCext_ VCC 47k
U115 __U115
C86 Ah GNDPWR 0.01m
XU117 VCC Net-_U101-_PE_ VCC Net-_U117-D1_ Net-_U117-D1_ Net-_U117-D3_ VCC GNDPWR Net-_U116-_PE_ _Vb Net-_U117-Q3_ Net-_U117-Q2_ Net-_U117-Q1_ Net-_U117-Q0_ VCC VCC NC-U117-0 NC-U117-1 NC-U117-2 74161
XU116 VCC Net-_U101-_PE_ GNDPWR GNDPWR GNDPWR GNDPWR VCC GNDPWR Net-_U116-_PE_ Net-_U116-CET_ Net-_U116-Q3_ Net-_U116-Q2_ Net-_U116-Q1_ Net-_U116-Q0_ VCC VCC NC-U116-0 NC-U116-1 NC-U116-2 74161
XU109 VCC Net-_U101-_PE_ GNDPWR GNDPWR GNDPWR GNDPWR VCC GNDPWR Net-_U104-_PE_ Net-_U104-TC_ Net-_U109-Q3_ Net-_U109-Q2_ Net-_U109-Q1_ Net-_U109-Q0_ VCC VCC NC-U109-0 NC-U109-1 NC-U109-2 74161
XU102 VCC 7MHz Net-_U102-D0_ Net-_U102-D1_ Net-_U102-D2_ Net-_U102-D3_ Net-_U102-CEP_ GNDPWR Net-_U101-_PE_ VCC Net-_U102-Q3_ Net-_U102-Q2_ Net-_U102-Q1_ Net-_U102-Q0_ VCC VCC NC-U102-0 NC-U102-1 NC-U102-2 74161
XU31 Net-_U20-CLR_ A26 7417
XU38 Net-_RN2H-R8.1_ VCC VCC Ak unconnected-_U38B-Q-Pad5_ Net-_U38B-Cext_ Net-_U38B-RCext_ Net-_U37A-_R_ Net-_U37A-_R_ 74123
XU29 Net-_U2-Pad3_ A20 7417
Cp25 GNDPWR VCC 100n
Cp38 GNDPWR VCC 100n
Cp39 GNDPWR VCC 100n
Cp22 GNDPWR VCC 100n
Cp18 GNDPWR VCC 100n
Cp23 GNDPWR VCC 100n
Cp1 GNDPWR VCC 100n
Cp15 GNDPWR VCC 100n
Cp10 GNDPWR VCC 100n
Cp34 GNDPWR VCC 100n
Cp31 GNDPWR VCC 100n
Cp33 GNDPWR VCC 100n
Cp13 GNDPWR VCC 100n
Cp14 GNDPWR VCC 100n
Cp19 GNDPWR VCC 100n
Cp32 GNDPWR VCC 100n
Cp30 GNDPWR VCC 100n
Cp40 GNDPWR VCC 100n
Cp12 GNDPWR VCC 100n
Cp37 GNDPWR VCC 100n
Cp17 GNDPWR VCC 100n
Cp26 GNDPWR VCC 100n
Cp28 GNDPWR VCC 100n
Cp24 GNDPWR VCC 100n
Cp11 GNDPWR VCC 100n
Cp20 GNDPWR VCC 100n
Cp29 GNDPWR VCC 100n
R21 VCC Net-_U121A-RCext_ 47k
XU121 Net-_U121A-A_ Net-_U121A-B_ Net-_U120A-Clr_ Net-_U121A-_Q_ Net-_U121A-A_ Net-_U121B-Cext_ Net-_U121B-RCext_ Net-_U121A-B_ Net-_U121A-B_ 74123
C34 Net-_U120A-RCext_ Net-_U120A-Cext_ 470m
R18 VCC Net-_U121B-RCext_ 47k
C32 Net-_U121B-RCext_ Net-_U121B-Cext_ 470m
C35 Net-_U121A-RCext_ Net-_U121A-Cext_ 470m
XU85 B21 Net-_U49A-Q_ unconnected-_U85-Pad3_ _L1-SIDE 7411
C31 Net-_U120B-RCext_ Net-_U120B-Cext_ 470m
R17 VCC Net-_U120B-RCext_ 47k
U40 U40.unbekannt
V1 VCC GNDPWR DC 1 
Cp27 GNDPWR VCC 100n
Cp35 GNDPWR VCC 100n
Cp36 GNDPWR VCC 100n
Cp21 GNDPWR VCC 100n
Cp2 GNDPWR VCC 100n
Cp5 GNDPWR VCC 100n
Cp4 GNDPWR VCC 100n
Cp6 GNDPWR VCC 100n
Cp8 GNDPWR VCC 100n
Cp16 GNDPWR VCC 100n
Cp7 GNDPWR VCC 100n
Cp9 GNDPWR VCC 100n
Cp3 GNDPWR VCC 100n
XU33 Net-_U33A-_R_ B9 Net-_U27B-Q_ VCC EXPLO._ST. _EXPLO._ST. 7474
XU37 Net-_U37A-_R_ VCC Net-_U20-_LOAD_ VCC B1 _COIN_IN 7474
XU89 Net-_U89-S_ GNDPWR VCC Net-_U89-Za_ GNDPWR Net-_U89-I1b_ Net-_U89-Zb_ GNDPWR Net-_U89-Zc_ Net-_U89-I1b_ GNDPWR Net-_U89-Zd_ Net-_U121A-B_ VCC VCC VCC NC-U89-0 NC-U89-1 NC-U89-2 NC-U89-3 NC-U89-4 NC-U89-5 NC-U89-6 74157
C4 Net-_U26-CV_ GNDPWR 0.1u
R4 Net-_U26-DIS_ Net-_U26-THR_ 12k
C5 Net-_U26-THR_ GNDPWR 47u
XU22 Net-_U22-Pad1_ Net-_U32D-Q_ Net-_U7-B3_ 7408
R5 Net-_R5-Pad1_ Net-_U26-DIS_ 3.3k
ARV1 Net-_R5-Pad1_ VCC unconnected-_RV1-Pad3_ __RV1
XU26 GNDPWR Net-_U26-THR_ Net-_U26-Q_ Net-_U26-R_ Net-_U26-CV_ Net-_U26-THR_ Net-_U26-DIS_ UA555
R998 Net-_D2-K_ A6 220
D2 VCC Net-_D2-K_ __D2
R22 VCC Net-_SW1-A_ 1k
SW1 __SW1
XU125 unconnected-_U125-Pad1_ unconnected-_U125-Pad2_ Net-_SW1-B_ Net-_U32A-Q_ 7411
XU32 Net-_U32A-_R_ Net-_RN2C-R3.1_ Net-_RN2C-R3.1_ Net-_U32A-Q_ Net-_RN2D-R4.1_ Net-_RN2E-R5.1_ Net-_U32B-Q_ 74279
XU12 Net-_U69-Za_ Net-_U10-Oa_b_ Net-_U25-UP_ 7400
XU21 74192
XU20 74192
C9 Net-_RN2E-R5.1_ GNDPWR 0.1u
C11 Net-_U32A-_R_ GNDPWR 470m
C37 Net-_U32C-_R_ GNDPWR 0.1m
R24 A32 Net-_U32C-_R_ 100
R23 VCC A32 560
C6 Net-_RN2D-R4.1_ GNDPWR 680p
C8 Net-_RN2C-R3.1_ GNDPWR 0.1u
RN2 Net-_RN2A-R1.1_ Net-_RN2B-R2.1_ 100
C12 Net-_RN2H-R8.1_ GNDPWR 0.01m
C14 Net-_RN2H-R8.1_ GNDPWR 47
SW5 __SW5
C13 Net-_RN2H-R8.1_ Net-_RN2H-R8.1_ 0.01m
R7 Net-_RN2H-R8.1_ VCC 100k
C19 Net-_U38A-RCext_ Net-_U38A-Cext_ 470m
R9 VCC Net-_U38A-RCext_ 47k
D1 Net-_D1-A_ Aj __D1
AE1 __AE1
C36 Net-_RN2G-R7.2_ GNDPWR 0.1m
XU50 Net-_U50A-_R_ VCC B2 unconnected-_U50A-_S-Pad4_ Net-_U50A-Q_ Net-_U50A-_Q_ 7474
QTR1 Net-_TR1-B_ A9 GNDPWR __TR1
XU90 VCC Net-_U101-_PE_ Net-_U89-Za_ Net-_U89-Zb_ Net-_U89-Zc_ Net-_U89-Zd_ VCC GNDPWR Net-_U90-_PE_ _Vb Net-_U90-Q3_ Net-_U90-Q2_ Net-_U90-Q1_ Net-_U90-Q0_ VCC VCC NC-U90-0 NC-U90-1 NC-U90-2 74161
R1 Net-_R1-Pad1_ Net-_TR1-B_ 560
R6 VCC A30 1k
C15 Net-_U38B-RCext_ Net-_U38B-Cext_ 0.1m
R8 VCC Net-_U38B-RCext_ 47k
XU55 Net-_C25-Pad1_ Net-_U55-Pad11_ B2 7432
L1 VCC A9 COIN METER
C25 Net-_C25-Pad1_ GNDPWR 1000p
R15 Net-_R15-Pad1_ Net-_C25-Pad1_ 220
XU79 74393
C41 A30 GNDPWR 470p
C27 Net-_C27-Pad1_ GNDPWR 1000p
R13 VCC Net-_U49A-RCext_ 47k
C24 Net-_U49A-RCext_ Net-_U49A-Cext_ 100m
XU49 B2 VCC VCC C1 _SPLAY_B Net-_U49B-Cext_ Net-_U49B-RCext_ CM CM 74123
R14 Net-_R14-Pad1_ Net-_C27-Pad1_ 220
XU27 unconnected-_U27A-_R-Pad1_ Net-_U27A-_S1_ Net-_U27A-_S1_ Net-_U27A-Q_ _HOME_POS.__G_ Net-_U27B-_S_ Net-_U27B-Q_ 74279
XU13 ACCE._D A12 7407
XU8 Vs/8 Net-_U7-Oa_b_ Net-_U15-DOWN_ 7400
U17 U17.unbekannt
U19 U19.unbekannt
U18 U18.unbekannt
XU28 unconnected-_U28-Pad1_ unconnected-_U28-Pad2_ Net-_U10-A1_ Net-_U10-A0_ 7410
XU2 Net-_U3-S0_ _SP._DOWN Net-_U2-Pad3_ 7408
XU43 CA PLAYER Net-_U15-QD_ Net-_U1A-A_ Net-_U43B-Q_ Net-_U43B-Cext_ Net-_U43B-RCext_ CM CM 74123
U16 __U16
C10 Net-_RN2B-R2.1_ GNDPWR 0.1u
XU6 Net-_U15-QD_ Net-_U6-Pad13_ 7404
XU23 EXPLO._ST. Net-_U27B-Q_ Net-_U4-_E_ 7432
XU1 Net-_U1A-A_ A8 Net-_U1A-Clr_ Net-_U1A-_Q_ Net-_U1B-Q_ Net-_U1B-Cext_ Net-_U1B-RCext_ Net-_U1A-A_ Net-_U1A-A_ 74123
XU14 ACCE._C ACCE._A NC-U14-0 ACCE._B unconnected-_U14-Pad5_ 7420
C7 Net-_RN2A-R1.1_ GNDPWR 0.1u
R11 VCC Net-_U43A-RCext_ 47k
C20 Net-_U43A-RCext_ Net-_U43A-Cext_ 10u
R10 VCC Net-_U43B-RCext_ 47k
XU9 74153
C2 Net-_U1A-RCext_ Net-_U1A-Cext_ 4.7m
R12 VCC Net-_U49B-RCext_ 47k
C21 Net-_U49B-RCext_ Net-_U49B-Cext_ 22m
C18 Net-_U43B-Cext_ Net-_U43B-RCext_ 15u
R2 VCC Net-_U1B-RCext_ 47k
C1 Net-_U1B-RCext_ Net-_U1B-Cext_ 4.7m
R3 VCC Net-_U1A-RCext_ 47k
XU67 B12 B12 Net-_U67B-2B_ B18 Net-_U67B-2D_ Net-_U5A-CP_ GNDPWR Net-_U67A-1Y_ B18 Net-_U67A-1D_ unconnected-_U67A-1X-Pad11_ unconnected-_U67A-1_X-Pad12_ VCC VCC NC-U67-0 NC-U67-1 NC-U67-2 7450
U11 __U11
U15 U15.unbekannt
U24 U24.unbekannt
U25 U25.unbekannt
U7 U7.unbekannt
U10 __U10
C16 Net-_U39A-CP_ GNDPWR 470p
U69 U69.unbekannt
XU60 Net-_U60-S_ B21 BX Net-_U60-Za_ B2 Vs/8 Net-_U60-Zb_ GNDPWR unconnected-_U60-Zc-Pad9_ unconnected-_U60-I1c-Pad10_ unconnected-_U60-I0c-Pad11_ unconnected-_U60-Zd-Pad12_ unconnected-_U60-I1d-Pad13_ unconnected-_U60-I0d-Pad14_ VCC VCC NC-U60-0 NC-U60-1 NC-U60-2 NC-U60-3 NC-U60-4 NC-U60-5 NC-U60-6 74157
C3 Net-_U19A-MR_ GNDPWR 470p
U5 __U5
XU4 Net-_U4-I2_ Net-_U4-I2_ Net-_U4-I0_ Net-_U4-I0_ Net-_U4-Z_ unconnected-_U4-_Z-Pad6_ Net-_U4-_E_ GNDPWR Net-_U10-B2_ Net-_U10-B1_ Net-_U10-B0_ Net-_U4-I6_ Net-_U4-I6_ Net-_U4-I4_ VCC VCC NC-U4-0 NC-U4-1 NC-U4-2 74151A
U42 U42.unbekannt
U36 __U36
U3 __U3
U35 U35.unbekannt
U41 __U41
U77 __U77
C17 Net-_U40A-MR_ GNDPWR 470p
.end
